interface design_out_intf (input clk);
	logic [9-1:0] x;
	logic [9-1:0] y;
	logic 		  valid;
endinterface 