interface design_in_intf (input clk);
	logic [7-1:0]a;
	logic [7-1:0]b;
	logic [7-1:0]c;
	logic 		 valid;	
	
endinterface 